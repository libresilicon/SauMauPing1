module testbench();
endmodule
